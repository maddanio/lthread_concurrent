module main

#flag -I @VMODROOT/src
#flag @VMODROOT/src/libcontext.o
#flag @VMODROOT/src/lthread.o
#flag @VMODROOT/src/lthread_cond.o
#flag @VMODROOT/src/lthread_socket.o
#flag @VMODROOT/src/lthread_poller.o

fn main() {
	println('Hello World!')
}
